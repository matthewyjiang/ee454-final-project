module cross_entropy_loss #(
    parameters
) (
    ports
);
    
endmodule